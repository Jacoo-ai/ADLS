`timescale 1ns / 1ps
module split2 #(
) (
    input logic data_in_valid,
    output logic data_in_ready,
    /* verilator lint_off UNOPTFLAT */
    output logic [1:0] data_out_valid,
    /* verilator lint_off UNOPTFLAT */
    input logic [1:0] data_out_ready
);
  // to make sure it can handshake correctly
  // only when in_valid && our_ready0 && out_ready1, handshake successfully
  // +-----------+-----------+------------+------------+------------+------------+
  // | in_valid  | outready0 | out_ready1 | out_valid0 | out_valid1 |  in_ready  |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         0 |         0 |          0 |          0 |          0 |          0 |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         0 |         0 |          1 |          0 |          0 |          0 |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         0 |         1 |          0 |          0 |          0 |          0 |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         0 |         1 |          1 |          0 |          0 |          1 |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         1 |         0 |          0 |          0 |          0 |          0 |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         1 |         0 |          1 |          1 |          0 |          0 |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         1 |         1 |          0 |          0 |          1 |          0 |
  // +-----------+-----------+------------+------------+------------+------------+
  // |         1 |         1 |          1 |          1 |          1 |          1 |
  // +-----------+-----------+------------+------------+------------+------------+
  always_comb begin
    data_out_valid[0] = data_in_valid && data_out_ready[1];
    data_out_valid[1] = data_in_valid && data_out_ready[0];
    data_in_ready     = data_out_ready[0] && data_out_ready[1];
  end
endmodule
